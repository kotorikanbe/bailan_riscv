module  Sixty_four_bit_multiplier 
    (
        input [63:0]      operator_1,
        input [63:0]      operator_2,
        output [63:0]     answer
    );

endmodule //Sixty_four_bit_multiplier